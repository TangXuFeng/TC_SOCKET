module dual_port_mem (
    input              clk,
    input              rst_n,

    // -------- Port 1: read + write --------
    input              write_1,
    input              read_1,
    input      [31:0]  address_1,
    input      [31:0]  write_data_1,
    output reg [31:0]  read_data_1,

    // -------- Port 2: read only --------
    input              read_2,
    input      [31:0]  address_2,
    output reg [31:0]  read_data_2
);

    // �ڴ��С������Ըĳ�����Ҫ�����
    localparam MEM_DEPTH = 1024;  // 1024 words = 4KB

    // 32-bit ��ȵ� RAM
    reg [31:0] mem [0:MEM_DEPTH-1];

    // ���ֽڵ�ַת��Ϊ word ��ַ
    wire [31:2] addr1_word = address_1[31:2];
    wire [31:2] addr2_word = address_2[31:2];

    // -----------------------------
    // Port 1: ͬ��д���첽��
    // -----------------------------
    always @(posedge clk) begin
        if (!rst_n) begin
            read_data_1 <= 32'b0;
        end else begin
            // д������ͬ����
            if (write_1) begin
                mem[addr1_word] <= write_data_1;
            end

            // ���������첽���Ĵ������
            if (read_1) begin
                read_data_1 <= mem[addr1_word];
            end
        end
    end

    // -----------------------------
    // Port 2: ֻ���˿�
    // -----------------------------
    always @(posedge clk) begin
        if (!rst_n) begin
            read_data_2 <= 32'b0;
        end else begin
            if (read_2) begin
                read_data_2 <= mem[addr2_word];
            end
        end
    end

endmodule

