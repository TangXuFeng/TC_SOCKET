module memory #(
 parameter SIZE = 20  // 2^20 bytes = 1MB
)(
 input              clk
 , input              rst_n

 , input              enable   // ѡ����
 , input              rw       // 0=��, 1=д
 , input      [31:0]  address
 , input      [31:0]  write_data
 , output reg wait_sig //�ȴ���,����д��æʱ����
 , output reg [31:0]  read_data
);

 // ---------------------------------------------------------
 // �ڴ����У�32bit ���
 // ���ֽ��� = 2^SIZE
 // �� word �� = 2^(SIZE-2)
 // ---------------------------------------------------------
 localparam WORDS = (1 << (SIZE - 2));

 reg [31:0] mem [0:WORDS-1];
 reg [4:0] wait_reg;

 // ---------------------------------------------------------
 // ��ַ���ֽ�Ѱַ����Ҫ���� 4 �õ� word index
 // ---------------------------------------------------------
 wire [31:0] word_index = address[31:2];

 // ---------------------------------------------------------
 // ͬ����д
 // ---------------------------------------------------------
 always @(posedge clk) begin
  if (!rst_n) begin
   read_data <= 32'b0;
   wait_reg<=5'b0;
  end else if (enable) begin
   //ģ���豸��æ,������16���ں󷵻�����
   //�ӳ��ڴ�
   wait_sig=1'b1;
   if(wait_reg == 5'b0)begin
    wait_reg<=wait_reg+5'b1;
   end else if(wait_reg == 5'b10000) begin
    wait_reg <= 5'b0;
    wait_sig= 1'b0;
   end
   if (rw == 1'b1) begin
    // д
    mem[word_index] <= write_data;
   end else begin
    // ��
    read_data <= mem[word_index];
   end
  end
 end

endmodule
