module riscv (
    input  clk
    ,input  rst_n
    ,input  in
    ,output pc
);

    // Core <-> dual_load_memory (I-port)
    wire [31:0] pc;
    wire [31:0] instruction;

    // Core <-> memory / dual_load_memory (D-port)
    wire [31:0] d_addr;
    wire [31:0] d_wdata;
    wire [31:0] d_rdata;
    wire        d_ren;
    wire        d_wen;

    // dual_load_memory outputs
    wire [31:0] dlm_rdata;
    wire        dlm_selected;

    // memory outputs
    wire [31:0] mem_rdata;
    wire        mem_selected;

    wire [31:0] external_interrupts; //�ⲿ�ж��ź�

    core #(
        .RST_PC_ADDRESS(32'h8000_0000)
    ) u_core (
        .clk            (clk)
        ,.rst_n          (rst_n)
        ,.pc             (pc)
        ,.instruction    (instruction)   // ���� dual_load_memory
        ,.external_interrupts   (external_interrupts)

        ,.address        (d_addr)
        ,.read_data      (d_rdata)       // ���� memory �� dual_load_memory
        ,.write_data     (d_wdata)
        ,.write_data_sig (d_wen)
    );

    dual_load_memory #(
        .MMIO_BASE_MEMORY(32'h8000_0000),
        .MMIO_MASK_MEMORY(32'hFFFF_FF00) //���볤�Ⱥ��ڴ��С�й�,2^8=256byte
    ) u_dual_load_memory (
        .clk        (clk),
        .rst_n      (rst_n),
        .pc         (pc),           // CPU ȡָ��ַ
        .instruction(instruction),  // ָ�����

        .address    (d_addr),       // CPU ���ݵ�ַ
        .read_data  (dlm_rdata),    // ���ݶ���
        .write_data (d_wdata),      // CPU д����
        .write_data_sig (d_wen),        // CPU д�ź�

        .selected   (dlm_selected)  // ��ַ����
    );

    memory #(
        .MMIO_BASE_MEMORY(32'h9000_0000),
        .MMIO_MASK_MEMORY(32'hFFFF_FF00) //���ڴ��ۺ�����������
    ) u_memory (
        .clk        (clk)
        ,.rst_n      (rst_n)

        ,.address    (d_addr)
        ,.read_data  (mem_rdata)
        ,.write_data (d_wdata)
        ,.write_data_sig         (d_wen)
        ,.selected   (mem_selected)
    );

    // ѡ����ĸ��豸��ȡ
    assign d_rdata = dlm_selected ? dlm_rdata 
                     :mem_selected ? mem_rdata
                     :32'b0;


endmodule
