module riscv (
    input  clk
    ,input  rst_n
    ,output done
);

// Core <-> dual_load_memory (I-port)
wire [31:0] pc;
wire [31:0] instruction;

// Core <-> memory / dual_load_memory (D-port)
wire [31:0] d_addr;
wire [31:0] d_wdata;
wire [31:0] d_rdata;
wire        d_ren;
wire        d_wen;

// dual_load_memory outputs
wire [31:0] dlm_rdata;
wire        dlm_selected;

// memory outputs
wire [31:0] mem_rdata;
wire        mem_selected;


    
core #(
    .RST_PC_ADDRESS(32'h0000_0000)
) u_core (
    .clk            (clk),
    .rst_n          (rst_n),

    .instruction    (instruction),   // ���� dual_load_memory
    .read_data      (d_rdata),       // ���� memory �� dual_load_memory

    .pc             (pc),
    .address        (d_addr),
    .write_data     (d_wdata),
    .read_data_sig  (d_ren),
    .write_data_sig (d_wen)
);
dual_load_memory #(
    .MMIO_BASE_MEMORY(32'h8000_0000),
    .MMIO_MASK_MEMORY(32'hFFFF_FF00) //���볤�Ⱥ��ڴ��С�й�,2^8=256byte
) u_dual_load_memory (
    .clk        (clk),
    .rst_n      (rst_n),

    .rw         (d_wen),        // CPU д�ź�
    .address    (d_addr),       // CPU ���ݵ�ַ
    .pc         (pc),           // CPU ȡָ��ַ
    .write_data (d_wdata),      // CPU д����

    .read_data  (dlm_rdata),    // ���ݶ���
    .instruction(instruction),  // ָ�����
    .selected   (dlm_selected)  // ��ַ����
);
memory #(
    .MMIO_BASE_MEMORY(32'h9000_0000),
    .MMIO_MASK_MEMORY(32'hFFFF_FF00) //���ڴ��ۺ�����������
) u_memory (
    .clk        (clk),
    .rst_n      (rst_n),

    .rw         (d_wen),
    .address    (d_addr),
    .write_data (d_wdata),

    .read_data  (mem_rdata),
    .selected   (mem_selected)
);

endmodule
