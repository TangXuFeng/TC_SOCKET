module alu #(
    parameter ENABLE_RV32M=0 //��ʿ,���Ҫ����Ӳ���˷�����?
)(
    input  [31:0] alu_a
    ,input  [31:0] alu_b
    ,input  [4:0]  alu_op

    ,output reg [31:0] alu_result
);


    parameter alu_add=  5'b00000;
    parameter alu_sll=  5'b00001;
    parameter alu_slt=  5'b00010;
    parameter alu_sltu= 5'b00011;
    parameter alu_xor=  5'b00100;
    parameter alu_srl=  5'b00101;
    parameter alu_or=   5'b00110;
    parameter alu_and=  5'b00111;
    
    parameter alu_sub=5'b01000;
    parameter alu_sra=  5'b01101;

    parameter alu_eq=5'b11000;

    parameter alu_mul=5'b10000;
    parameter alu_mulh=5'b10001;
    parameter alu_mulhsu=5'b10010;
    parameter alu_mulhu=5'b10011;
    parameter alu_div=5'b10100;
    parameter alu_divu=5'b10101;
    parameter alu_rem=5'b10110;
    parameter alu_remu=5'b10111;

    reg [63:0] tmp;
    always @(*)begin
        alu_result = 32'b0;
        tmp = 64'b0;

        if(alu_op==alu_add || alu_op==alu_sub)alu_result = alu_a + alu_op[3]?-alu_b:alu_b;
        if(alu_op[4:3] == 2'b00)begin
            case(alu_op[2:0])
                3'b001:alu_result = alu_a << alu_b[4:0];
                3'b010:alu_result = $signed(alu_a) < $signed(alu_b)?32'b1:32'b0; 
                3'b011:alu_result = alu_a < alu_b ? 32'b1:32'b0;
                3'b100:alu_result = alu_a ^ alu_b;
                3'b110:alu_result = alu_a | alu_b;
                3'b111:alu_result = alu_a & alu_b;
            endcase
        end
        if(alu_op==alu_sra) alu_result =  $signed(alu_a) >>> alu_b[4:0]; 
        if(alu_op==alu_eq)  alu_result = alu_a == alu_b ? 32'b1:32'b0;


        // �˷����ͳ�����������Ū���жϴ�������ڳ�����
        //generate
            //TCʵ����Ϊ�˽�Լ�����˷����ͳ�����
            //���������ж��Ƿ��Ǹ���
            //Ȼ��ȡ����ֵ(����Ǹ���,��ȡ��,�������)
            //�����,������������ж��Ƿ���Ҫ�ٴ�ȡ��
            //�����˳��������Ϊ����,��Ҫȡ���ָ������ȷ��
            //�����˳�����,�����˳��������Ϊ��,����ȡ��
            if(ENABLE_RV32M)begin
                if(alu_op[4:3]==2'b10)begin
                    case(alu_op[2:0])
                        3'b000,3'b001:tmp = (alu_a*alu_b);
                        3'b010:tmp = $signed(alu_a) * alu_b;
                        3'b011:tmp = $signed(alu_a) * $signed(alu_b);

                        3'b100:tmp = (alu_b == 0) ? 32'hFFFFFFFF : $signed(alu_a) / $signed(alu_b);
                        3'b101:tmp = (alu_b == 0) ? 32'hFFFFFFFF : alu_a / alu_b;
                        3'b110:tmp = (alu_b == 0) ? alu_a : $signed(alu_a) % $signed(alu_b);
                        3'b111:tmp = (alu_b == 0) ? alu_a : alu_a % alu_b;
                    endcase
                    if(alu_op[2:0]==3'b0 || alu_op[2:1]==3'b10)alu_result=tmp[31:0];
                    else alu_result=tmp[63:0];
                end
            end else begin
                //�����жϴ���
            end
        //endgenerate


    end
endmodule

