module alu #(
    parameter ENABLE_RV32M=0 //��ʿ,���Ҫ����Ӳ���˷�����?
)(
    input  [31:0] alu_a
    ,input  [31:0] alu_b
    ,input  [5:0]  alu_op

    ,output reg [31:0] alu_result
);
    //alu_op:
    //�����ж�1'b1,funct7[0]  ,funct7[5],funct3[2:0]


    parameter alu_add=  5'b00000;
    parameter alu_sll=  5'b00001;
    parameter alu_xor=  5'b00100;
    parameter alu_srl=  5'b00101;
    parameter alu_or=   5'b00110;
    parameter alu_and=  5'b00111;

    parameter alu_sub=5'b01000;
    parameter alu_sra=  5'b01101;


    parameter alu_mul=5'b10000;
    parameter alu_mulh=5'b10001;
    parameter alu_mulhsu=5'b10010;
    parameter alu_mulhu=5'b10011;
    parameter alu_div=5'b10100;
    parameter alu_divu=5'b10101;
    parameter alu_rem=5'b10110;
    parameter alu_remu=5'b10111;

    reg [63:0] tmp;

    wire eq  = alu_a == alu_b;
    wire lt  = $signed(alu_a) < $signed(alu_b);
    wire ltu = alu_a < alu_b;

    always @(*)begin
        alu_result = 32'b0;
        tmp = 64'b0;
        if(alu_op[5]==1'b1)begin

            //beq  000 a=b
            //bne  001 a!=b 
            //bge  101 a>=b signed
            //bgeu 111 a>=b unsigned
            //blt  100 a<b  signed
            //bltu 110 a<b  unsigned           
            alu_result = (alu_op[0]^(alu_op[2]?(alu_op[1]?lt:ltu):eq))?32'b1:32'b0;

        end else begin
            if(alu_op[4] == 1'b0)begin
                case(alu_op[2:0])
                    3'b000:alu_result = alu_a + (alu_op[3]?-alu_b +1:alu_b); //add sub
                    3'b001:alu_result = alu_a << alu_b[4:0]; //sll
                    3'b010:alu_result = lt?32'b1:32'b0; 
                    3'b011:alu_result = ltu ? 32'b1:32'b0;
                    3'b100:alu_result = alu_a ^ alu_b;
                    3'b101:alu_result = alu_op[3]?$signed(alu_a) >>> alu_b[4:0]:alu_a >> alu_b[4:0];
                    3'b110:alu_result = alu_a | alu_b;
                    3'b111:alu_result = alu_a & alu_b;
                endcase
            end


            // �˷����ͳ�����������Ū���жϴ�������ڳ�����
            //generate
            //TCʵ����Ϊ�˽�Լ�����˷����ͳ�����
            //���������ж��Ƿ��Ǹ���
            //Ȼ��ȡ����ֵ(����Ǹ���,��ȡ��,�������)
            //�����,������������ж��Ƿ���Ҫ�ٴ�ȡ��
            //�����˳��������Ϊ����,��Ҫȡ���ָ������ȷ��
            //�����˳�����,�����˳��������Ϊ��,����ȡ��
            if(ENABLE_RV32M)begin
                if(alu_op[4:3]==2'b10)begin
                    case(alu_op[2:0])
                        3'b000,3'b001:tmp = (alu_a*alu_b);
                        3'b010:tmp = $signed(alu_a) * alu_b;
                        3'b011:tmp = $signed(alu_a) * $signed(alu_b);

                        3'b100:tmp = (alu_b == 0) ? 32'hFFFFFFFF : $signed(alu_a) / $signed(alu_b);
                        3'b101:tmp = (alu_b == 0) ? 32'hFFFFFFFF : alu_a / alu_b;
                        3'b110:tmp = (alu_b == 0) ? alu_a : $signed(alu_a) % $signed(alu_b);
                        3'b111:tmp = (alu_b == 0) ? alu_a : alu_a % alu_b;
                    endcase
                    if(alu_op[2:0]==3'b0 || alu_op[2:1]==3'b10)alu_result=tmp[31:0];
                    else alu_result=tmp[63:0];
                end
            end else begin
                //�����жϴ���
            end
            //endgenerate
        end
    end
endmodule

