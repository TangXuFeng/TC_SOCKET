//˫�����ڴ�
module dual_load_memory #(
    parameter MMIO_BASE_MEMORY = 32'h80000000 //����ַ
    ,parameter MMIO_MASK_MEMORY = 32'hFFFFFF00 //����
)(
    input               clk
    ,input              rst_n

    ,input              rw       // 0=��, 1=д
    ,input      [31:0]  address
    ,input      [31:0]  pc
    ,input      [31:0]  write_data

    ,output     [31:0]  read_data // �첽��
    ,output     [31:0]  instruction
    ,output             selected //ѡ���ź�
);
    //�����ڴ��С
    localparam MEM_SIZE = (~MMIO_MASK_MEMORY)>>2 +1;
    reg [31:0] mem [0:MEM_SIZE];
    wire selected_instruction= (address & MMIO_MASK_MEMORY)==MMIO_BASE_MEMORY;
    assign selected = (address & MMIO_MASK_MEMORY)==MMIO_BASE_MEMORY;

    assign instruction=(selected_instruction && pc[1:0]==0 ) ? mem[address[31:2]] : 32'b0;

    //��ȡ,���ҵ�λ��ַ�������0
    assign read_data = (selected && rw == 1'b0 && address[1:0]==0 ) ? mem[address[31:2]] : 32'b0;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            //��װ������
            mem[0]=32'b0;
        end else if (selected &&rw == 1'b1 && address[1:0] == 2'b00) begin
            mem[address[31:2]] <= write_data;
        end
    end

endmodule
