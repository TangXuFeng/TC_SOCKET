module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_1[7:0]), .en(wire_64), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_95), .in(arch_input_value), .out(wire_56));
  TC_Register # (.UUID(64'd3567277318659926168 ^ UUID), .BIT_WIDTH(64'd8)) Register8_2 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_74), .in(wire_1[7:0]), .out(wire_19));
  TC_Register # (.UUID(64'd4314171501159748010 ^ UUID), .BIT_WIDTH(64'd8)) Register8_3 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_12), .in(wire_1[7:0]), .out(wire_82));
  TC_Register # (.UUID(64'd4600363545443072287 ^ UUID), .BIT_WIDTH(64'd8)) Register8_4 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_54), .in(wire_1[7:0]), .out(wire_109));
  TC_Register # (.UUID(64'd730748584646115835 ^ UUID), .BIT_WIDTH(64'd8)) Register8_5 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_90), .in(wire_1[7:0]), .out(wire_65));
  TC_Splitter8 # (.UUID(64'd1498371318102751634 ^ UUID)) Splitter8_6 (.in(wire_22[7:0]), .out0(wire_26), .out1(wire_51), .out2(wire_80), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3337292616224932375 ^ UUID)) Decoder3_7 (.dis(wire_10), .sel0(wire_26), .sel1(wire_51), .sel2(wire_80), .out0(wire_113), .out1(wire_58), .out2(wire_66), .out3(wire_103), .out4(wire_5), .out5(wire_104), .out6(wire_37), .out7(wire_27));
  TC_Switch # (.UUID(64'd1917227579263597525 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_113), .in(wire_19), .out(wire_14_0));
  TC_Switch # (.UUID(64'd4606595889790715338 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_99), .in(wire_19), .out(wire_13_1));
  TC_Switch # (.UUID(64'd2755432556508539602 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_58), .in(wire_82), .out(wire_14_1));
  TC_Switch # (.UUID(64'd1283073392276043494 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_108), .in(wire_82), .out(wire_13_2));
  TC_Switch # (.UUID(64'd1028020839011630262 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_66), .in(wire_109), .out(wire_14_2));
  TC_Switch # (.UUID(64'd1679043610028313863 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_49), .in(wire_109), .out(wire_13_3));
  TC_Switch # (.UUID(64'd1594805671157965134 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_103), .in(wire_55), .out(wire_14_3));
  TC_Switch # (.UUID(64'd218360417323196330 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_45), .in(wire_55), .out(wire_13_4));
  TC_Switch # (.UUID(64'd3091015626988790686 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_5), .in(wire_65), .out(wire_14_5));
  TC_Switch # (.UUID(64'd3560473234436325609 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_33), .in(wire_65), .out(wire_13_5));
  TC_Switch # (.UUID(64'd3904266495292750520 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_104), .in(wire_79), .out(wire_14_6));
  TC_Switch # (.UUID(64'd2412792690051011461 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_114), .in(wire_79), .out(wire_13_6));
  TC_Or # (.UUID(64'd524826494083966693 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_83), .in1(wire_27), .out(wire_95));
  TC_Switch # (.UUID(64'd997672195784530257 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_37), .in(wire_28), .out(wire_14_7));
  TC_Switch # (.UUID(64'd376390880793986874 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_62), .in(wire_28), .out(wire_13_7));
  TC_Switch # (.UUID(64'd1523442411670562667 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_27), .in(wire_56), .out(wire_14_8));
  TC_Switch # (.UUID(64'd234999404583407884 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_83), .in(wire_56), .out(wire_13_8));
  TC_Splitter8 # (.UUID(64'd4424477377516370233 ^ UUID)) Splitter8_25 (.in(wire_44[7:0]), .out0(wire_50), .out1(wire_35), .out2(wire_106), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2689837594562073296 ^ UUID)) Decoder3_26 (.dis(wire_40), .sel0(wire_50), .sel1(wire_35), .sel2(wire_106), .out0(wire_99), .out1(wire_108), .out2(wire_49), .out3(wire_45), .out4(wire_33), .out5(wire_114), .out6(wire_62), .out7(wire_83));
  TC_Splitter8 # (.UUID(64'd240125590333452382 ^ UUID)) Splitter8_27 (.in(wire_4[7:0]), .out0(wire_53), .out1(wire_17), .out2(wire_124), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3641953999819191224 ^ UUID)) Decoder3_28 (.dis(wire_60), .sel0(wire_53), .sel1(wire_17), .sel2(wire_124), .out0(wire_74), .out1(wire_12), .out2(wire_54), .out3(wire_23), .out4(wire_90), .out5(wire_46), .out6(wire_111), .out7(wire_64));
  TC_Constant # (.UUID(64'd33792831588053931 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_29 (.out(wire_34));
  TC_Splitter8 # (.UUID(64'd3880695259190352202 ^ UUID)) Splitter8_30 (.in(wire_0[7:0]), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(wire_40), .out7(wire_10));
  TC_Switch # (.UUID(64'd4170108392612781585 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_10), .in(wire_22[7:0]), .out(wire_14_4));
  TC_Switch # (.UUID(64'd2160572697214472976 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_40), .in(wire_44[7:0]), .out(wire_13_0));
  TC_Mux # (.UUID(64'd321366353718168891 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_33 (.sel(wire_16), .in0(wire_1[7:0]), .in1(wire_4[7:0]), .out(wire_88));
  TC_Or # (.UUID(64'd3698707902444612499 ^ UUID), .BIT_WIDTH(64'd1)) Or_34 (.in0(wire_111), .in1(wire_16), .out(wire_29));
  TC_Program # (.UUID(64'd3443569880668636320 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_2FCA048FC87D04A0.w8.bin"), .ARG_SIG("Program_2FCA048FC87D04A0=%s")) Program_35 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_28 }), .out0(wire_0), .out1(wire_22), .out2(wire_44), .out3(wire_4));
  TC_Register # (.UUID(64'd386228554135477644 ^ UUID), .BIT_WIDTH(64'd8)) Register8_36 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_46), .in(wire_1[7:0]), .out(wire_79));
  TC_Register # (.UUID(64'd4342942410494833631 ^ UUID), .BIT_WIDTH(64'd8)) Register8_37 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_23), .in(wire_1[7:0]), .out(wire_55));
  TC_Splitter8 # (.UUID(64'd135032747788271218 ^ UUID)) Splitter8_38 (.in(wire_0[7:0]), .out0(), .out1(), .out2(), .out3(wire_89), .out4(wire_73), .out5(wire_39), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd4434827245328719037 ^ UUID)) Decoder3_39 (.dis(1'd0), .sel0(wire_89), .sel1(wire_73), .sel2(wire_39), .out0(wire_100), .out1(wire_72), .out2(wire_107), .out3(wire_92), .out4(wire_117), .out5(wire_25), .out6(wire_42), .out7(wire_63));
  TC_Maker8 # (.UUID(64'd1666200326811008964 ^ UUID)) Maker8_40 (.in0(wire_100), .in1(wire_72), .in2(wire_107), .in3(wire_92), .in4(wire_117), .in5(wire_25), .in6(wire_42), .in7(wire_63), .out(wire_97));
  TC_Not # (.UUID(64'd2777290053930372847 ^ UUID), .BIT_WIDTH(64'd8)) Not8_41 (.in(wire_97), .out(wire_36));
  TC_Splitter8 # (.UUID(64'd1067884220173821292 ^ UUID)) Splitter8_42 (.in(wire_36), .out0(wire_52), .out1(), .out2(), .out3(), .out4(wire_6), .out5(), .out6(), .out7(wire_93));
  TC_Splitter8 # (.UUID(64'd4567134934692615408 ^ UUID)) Splitter8_43 (.in(wire_0[7:0]), .out0(wire_59), .out1(wire_126), .out2(wire_98), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd1694196926993949689 ^ UUID)) Decoder3_44 (.dis(wire_93), .sel0(wire_59), .sel1(wire_126), .sel2(wire_98), .out0(), .out1(), .out2(), .out3(), .out4(wire_57), .out5(wire_91), .out6(wire_110), .out7(wire_61));
  TC_Nor # (.UUID(64'd4330657655357727171 ^ UUID), .BIT_WIDTH(64'd1)) Nor_45 (.in0(wire_91), .in1(wire_61), .out(wire_43));
  TC_Switch # (.UUID(64'd1003947045976264357 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_46 (.en(wire_43), .in(wire_52), .out(wire_60));
  TC_Counter # (.UUID(64'd3697303885325073163 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_47 (.clk(clk), .rst(rst), .save(wire_29), .in(wire_88), .out(wire_28));
  ZXE6ZXA0ZX88z_2 # (.UUID(64'd1958025861551982969 ^ UUID)) ZXE6ZXA0ZX88z_2_48 (.clk(clk), .rst(rst), .POP(wire_61), .PUSH(wire_110), .VALUE(wire_13), .OUTPUT(wire_1_8[7:0]));
  TC_Ram # (.UUID(64'd1129193633547332749 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_49 (.clk(clk), .rst(rst), .load(wire_91), .save(wire_57), .address({{24{1'b0}}, wire_14 }), .in0({{56{1'b0}}, wire_13 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_1_7), .out1(), .out2(), .out3());
  TC_Buffer # (.UUID(64'd3947718059578401630 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_50 (.in(wire_0[7:0]), .out(wire_120));
  TC_Buffer # (.UUID(64'd1704804697455945226 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_51 (.in(wire_14), .out(wire_47));
  TC_Buffer # (.UUID(64'd267809227722467906 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_52 (.in(wire_13), .out(wire_15));
  TC_Equal # (.UUID(64'd2232146239500284594 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_53 (.in0(wire_47), .in1(wire_15), .out(wire_24));
  TC_Splitter8 # (.UUID(64'd2849055587936809322 ^ UUID)) Splitter8_54 (.in(wire_120), .out0(wire_121), .out1(wire_18), .out2(wire_112), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3059271986324868397 ^ UUID)) Decoder3_55 (.dis(wire_123), .sel0(wire_121), .sel1(wire_18), .sel2(wire_112), .out0(wire_30), .out1(wire_32), .out2(wire_105), .out3(wire_86), .out4(wire_41), .out5(wire_75), .out6(), .out7());
  TC_Switch # (.UUID(64'd1448046988067494572 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_56 (.en(wire_30), .in(wire_24), .out(wire_16_5));
  TC_Not # (.UUID(64'd2613994107786124569 ^ UUID), .BIT_WIDTH(64'd1)) Not_57 (.in(wire_24), .out(wire_67));
  TC_Switch # (.UUID(64'd4291545752474881129 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_58 (.en(wire_32), .in(wire_67), .out(wire_16_4));
  TC_LessU # (.UUID(64'd4492936371535056576 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_59 (.in0(wire_47), .in1(wire_15), .out(wire_38));
  TC_Switch # (.UUID(64'd3204093226559410080 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_60 (.en(wire_105), .in(wire_38), .out(wire_16_3));
  TC_Or # (.UUID(64'd49567376829383419 ^ UUID), .BIT_WIDTH(64'd1)) Or_61 (.in0(wire_38), .in1(wire_24), .out(wire_48));
  TC_Switch # (.UUID(64'd2601095734074638618 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_62 (.en(wire_86), .in(wire_48), .out(wire_16_2));
  TC_Not # (.UUID(64'd1125903052844312452 ^ UUID), .BIT_WIDTH(64'd1)) Not_63 (.in(wire_24), .out(wire_102));
  TC_Not # (.UUID(64'd4584840909470784956 ^ UUID), .BIT_WIDTH(64'd1)) Not_64 (.in(wire_38), .out(wire_71));
  TC_And # (.UUID(64'd1416909615970935125 ^ UUID), .BIT_WIDTH(64'd1)) And_65 (.in0(wire_102), .in1(wire_71), .out(wire_96));
  TC_Switch # (.UUID(64'd1339841755482262318 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_66 (.en(wire_41), .in(wire_96), .out(wire_16_1));
  TC_Or # (.UUID(64'd2888452720716452071 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_24), .in1(wire_84), .out(wire_125));
  TC_Not # (.UUID(64'd1724070206610901975 ^ UUID), .BIT_WIDTH(64'd1)) Not_68 (.in(wire_38), .out(wire_84));
  TC_Switch # (.UUID(64'd3091203752929709012 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_69 (.en(wire_75), .in(wire_125), .out(wire_16_0));
  TC_Buffer # (.UUID(64'd2644856339883139859 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_70 (.in(wire_16), .out());
  TC_Buffer # (.UUID(64'd2924922131119042023 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_71 (.in(wire_6), .out(wire_123));
  TC_Buffer # (.UUID(64'd170079748537936221 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_72 (.in(wire_14), .out(wire_3));
  TC_Buffer # (.UUID(64'd2208771414383649028 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_73 (.in(wire_13), .out(wire_2));
  TC_Buffer # (.UUID(64'd3451990466605623828 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_74 (.in(wire_0[7:0]), .out(wire_94));
  TC_Add # (.UUID(64'd1401776941361291601 ^ UUID), .BIT_WIDTH(64'd8)) Add8_75 (.in0(wire_3), .in1(wire_8), .ci(wire_69), .out(wire_101), .co());
  TC_Splitter8 # (.UUID(64'd362369203052203362 ^ UUID)) Splitter8_76 (.in(wire_94), .out0(wire_69), .out1(wire_20), .out2(wire_122), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Mux # (.UUID(64'd3469026213967727577 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_77 (.sel(wire_69), .in0(wire_2), .in1(wire_70), .out(wire_8));
  TC_Not # (.UUID(64'd2498644868945124409 ^ UUID), .BIT_WIDTH(64'd8)) Not8_78 (.in(wire_2), .out(wire_70));
  TC_Switch # (.UUID(64'd545664435932097951 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_79 (.en(wire_81), .in(wire_101), .out(wire_1_5[7:0]));
  TC_And # (.UUID(64'd1249309791502122121 ^ UUID), .BIT_WIDTH(64'd8)) And8_80 (.in0(wire_3), .in1(wire_2), .out(wire_85));
  TC_Or # (.UUID(64'd206422988164098941 ^ UUID), .BIT_WIDTH(64'd8)) Or8_81 (.in0(wire_3), .in1(wire_2), .out(wire_87));
  TC_Not # (.UUID(64'd2239308705472345375 ^ UUID), .BIT_WIDTH(64'd8)) Not8_82 (.in(wire_3), .out(wire_11));
  TC_Xor # (.UUID(64'd4006105807823375779 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_83 (.in0(wire_3), .in1(wire_2), .out(wire_116));
  TC_Switch # (.UUID(64'd3756800535143481882 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_84 (.en(wire_76), .in(wire_85), .out(wire_1_3[7:0]));
  TC_Switch # (.UUID(64'd1039941532573398485 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_85 (.en(wire_118), .in(wire_87), .out(wire_1_0[7:0]));
  TC_Switch # (.UUID(64'd363584717263902295 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_86 (.en(wire_7), .in(wire_11), .out(wire_1_1[7:0]));
  TC_Switch # (.UUID(64'd384703047578586851 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_87 (.en(wire_21), .in(wire_116), .out(wire_1_2[7:0]));
  TC_Decoder3 # (.UUID(64'd550532555031177802 ^ UUID)) Decoder3_88 (.dis(wire_77), .sel0(wire_69), .sel1(wire_20), .sel2(wire_122), .out0(wire_31), .out1(wire_78), .out2(wire_76), .out3(wire_118), .out4(wire_7), .out5(wire_21), .out6(wire_119), .out7(wire_115));
  TC_Or # (.UUID(64'd3540251693030169431 ^ UUID), .BIT_WIDTH(64'd1)) Or_89 (.in0(wire_31), .in1(wire_78), .out(wire_81));
  TC_Buffer # (.UUID(64'd3619107362250460489 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_90 (.in(wire_52), .out(wire_77));
  TC_Buffer # (.UUID(64'd1031596948683568636 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_91 (.in(wire_1[7:0]), .out());
  TC_Shl # (.UUID(64'd3329634151053019757 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_92 (.in(wire_3), .shift(wire_2), .out(wire_9));
  TC_Shr # (.UUID(64'd2757397292058891751 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_93 (.in(wire_3), .shift(wire_2), .out(wire_68));
  TC_Switch # (.UUID(64'd4185839264255496959 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_94 (.en(wire_119), .in(wire_9), .out(wire_1_4[7:0]));
  TC_Switch # (.UUID(64'd2438550331752004072 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_95 (.en(wire_115), .in(wire_68), .out(wire_1_6[7:0]));

  wire [63:0] wire_0;
  wire [63:0] wire_1;
  wire [63:0] wire_1_0;
  wire [63:0] wire_1_1;
  wire [63:0] wire_1_2;
  wire [63:0] wire_1_3;
  wire [63:0] wire_1_4;
  wire [63:0] wire_1_5;
  wire [63:0] wire_1_6;
  wire [63:0] wire_1_7;
  wire [63:0] wire_1_8;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [63:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_13_0;
  wire [7:0] wire_13_1;
  wire [7:0] wire_13_2;
  wire [7:0] wire_13_3;
  wire [7:0] wire_13_4;
  wire [7:0] wire_13_5;
  wire [7:0] wire_13_6;
  wire [7:0] wire_13_7;
  wire [7:0] wire_13_8;
  assign wire_13 = wire_13_0|wire_13_1|wire_13_2|wire_13_3|wire_13_4|wire_13_5|wire_13_6|wire_13_7|wire_13_8;
  wire [7:0] wire_14;
  wire [7:0] wire_14_0;
  wire [7:0] wire_14_1;
  wire [7:0] wire_14_2;
  wire [7:0] wire_14_3;
  wire [7:0] wire_14_4;
  wire [7:0] wire_14_5;
  wire [7:0] wire_14_6;
  wire [7:0] wire_14_7;
  wire [7:0] wire_14_8;
  assign wire_14 = wire_14_0|wire_14_1|wire_14_2|wire_14_3|wire_14_4|wire_14_5|wire_14_6|wire_14_7|wire_14_8;
  wire [7:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_16_0;
  wire [0:0] wire_16_1;
  wire [0:0] wire_16_2;
  wire [0:0] wire_16_3;
  wire [0:0] wire_16_4;
  wire [0:0] wire_16_5;
  assign wire_16 = wire_16_0|wire_16_1|wire_16_2|wire_16_3|wire_16_4|wire_16_5;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [63:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [63:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [7:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [7:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  assign arch_output_enable = wire_64;
  wire [7:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  wire [0:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [7:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [7:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [7:0] wire_85;
  wire [0:0] wire_86;
  wire [7:0] wire_87;
  wire [7:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [7:0] wire_94;
  wire [0:0] wire_95;
  assign arch_input_enable = wire_95;
  wire [0:0] wire_96;
  wire [7:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [7:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [7:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [0:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [7:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [0:0] wire_126;

endmodule
