module memory #(
    parameter SIZE = 20  // 2^20 bytes = 1MB
)(
    input              clk,
    input              rst_n,

    input              enable,   // ѡ����
    input              rw,       // 0=��, 1=д
    input      [31:0]  address,
    input      [31:0]  write_data,

    output reg         wait_sig, // �ȴ���
    output     [31:0]  read_data, // �첽��
    output reg         instruction_address_misaligned
);

    // ---------------------------------------------------------
    // �ڴ����У�32bit ���
    // ���ֽ��� = 2^SIZE
    // �� word �� = 2^(SIZE-2)
    // ---------------------------------------------------------
    localparam WORDS = (1 << (SIZE - 2));

    reg [31:0] mem [0:WORDS-1];
    reg [4:0] wait_reg;

    // ---------------------------------------------------------
    // ��ַ���ֽ�Ѱַ����Ҫ���� 4 �õ� word index
    // ---------------------------------------------------------
    wire [31:0] word_index = address[31:2];

    // ---------------------------------------------------------
    //  �첽��������߼�ֱ�����
    // ---------------------------------------------------------
    assign read_data = (enable && rw == 1'b0) ? mem[word_index] : 32'b0;

    // ---------------------------------------------------------
    //  ͬ��д + �쳣��� + wait_sig ģ���ӳ�
    // ---------------------------------------------------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            instruction_address_misaligned <= 1'b0;
            wait_sig <= 1'b0;
            wait_reg <= 5'b0;
        end else begin

            // Ĭ�����쳣
            instruction_address_misaligned <= 1'b0;

            if (enable) begin

                // -------------------------------
                // ��ַδ�����쳣
                // -------------------------------
                if (address[1:0] != 2'b00) begin
                    instruction_address_misaligned <= 1'b1;
                end

                // -------------------------------
                // ģ���豸�ӳ٣�16 ����
                // -------------------------------
                if (wait_reg == 5'b0) begin
                    wait_sig <= 1'b1;
                    wait_reg <= wait_reg + 1'b1;
                end else if (wait_reg == 5'b10000) begin
                    wait_sig <= 1'b0;
                    wait_reg <= 5'b0;
                end else begin
                    wait_reg <= wait_reg + 1'b1;
                end

                // -------------------------------
                //  ͬ��д
                // -------------------------------
                if (rw == 1'b1 && address[1:0] == 2'b00) begin
                    mem[word_index] <= write_data;
                end
            end else begin
                wait_sig <= 1'b0;
                wait_reg <= 5'b0;
            end
        end
    end

endmodule
