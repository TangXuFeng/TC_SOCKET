module memory #(
    parameter MMIO_BASE_MEMORY = 32'h80000000 //����ַ
    ,parameter MMIO_MASK_MEMORY = 32'hFFF00000 //���� 20bit = 1MB
)(
    input               clk
    ,input              rst_n

    ,input              rw       // 0=��, 1=д
    ,input      [31:0]  address
    ,input      [31:0]  write_data

    ,output     [31:0]  read_data // �첽��
    ,output             interruped_0 //0���쳣,�ڴ治����:
    ,output             selected //ѡ���ź�
    ,output     [1:0]   cache_allow //֪ͨcache���ܱ�����,bit0��д����,bit1�Ƕ�����
);
    //�����ڴ��С
    localparam MEM_SIZE = (~MMIO_MASK_MEMORY)+1;
    reg [31:0] mem [MEM_SIZE:0];

    assign selected = (address & MMIO_MASK_MEMORY)==MMIO_BASE_MEMORY;
    assign interruped_0 = address[1:0] !=2'b0;
    assign cache_allow = selected? 2'b11:2'b11; //���Ա�����

    //��ȡ,���ҵ�λ��ַ�������0
    assign read_data = (selected && rw == 1'b0 && address[1:0]==0 ) ? mem[address[31:2]] : 32'b0;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            //��װ������
            mem[0]=32'b0;
        end else if (selected &&rw == 1'b1 && address[1:0] == 2'b00) begin
            mem[address[31:2]] <= write_data;
        end
    end

endmodule
