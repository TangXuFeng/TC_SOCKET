module memory_controller (
    input         clk
    , input         rst_n

    // ���� core �ķô�����
    , input         mem_read
    , input         mem_write
    , input  [31:0] mem_address
    , input  [31:0] mem_write_data
    , input  [2:0]  mem_size        // 0=1B, 1=2B, 3=4B

    // ���ظ� core
    , output reg [31:0] mem_read_data
    , output reg        mem_wait    // 1=æ��core ����ȴ�

    // ----------- ���ӵ� memory��dual_port_mem��-----------
    // ͨ��1����д
    , output reg        ch1_read
    , output reg        ch1_write
    , output reg [31:0] ch1_addr
    , output reg [31:0] ch1_wdata
    , input      [31:0] ch1_rdata

    // ͨ��2�����صڶ��� word ���ж�д
    , output reg        ch2_read
    , output reg [31:0] ch2_addr
    , input      [31:0] ch2_rdata
);

    // -------------------------
    // �����ֽ������Ƿ�� word
    // -------------------------
    wire [1:0] offset    = mem_address[1:0];

    wire [2:0] size_bytes =
        (mem_size == 3'd0) ? 3'd1 :
        (mem_size == 3'd1) ? 3'd2 :
        (mem_size == 3'd3) ? 3'd4 : 3'd4;  // ����ֵ�� 4 �ֽڴ���

    wire       cross_word = (offset + size_bytes) > 3'd4;

    wire [31:0] base_addr = {mem_address[31:2], 2'b00};
    wire [31:0] next_addr = base_addr + 32'd4;

    // -------------------------
    // FSM ״̬
    // -------------------------
    localparam S_IDLE        = 2'd0;
    localparam S_PHASE1      = 2'd1;  // �ѷ����һ�η��ʣ�������
    localparam S_PHASE2      = 2'd2;  // ���õ���һ word������ڶ� word

    reg [1:0] state;

    // �����һ�ζ����� 32bit
    reg [31:0] buffer;

    // ��¼��ǰ�����Ƕ�����д
    reg op_read;
    reg op_write;
    reg [31:0] latched_addr;
    reg [2:0]  latched_size;
    reg [31:0] latched_wdata;

    // -------------------------
    // ��ʱ���߼�
    // -------------------------
    always @(posedge clk) begin
        if (!rst_n) begin
            state        <= S_IDLE;
            mem_wait     <= 1'b0;

            ch1_read     <= 1'b0;
            ch1_write    <= 1'b0;
            ch2_read     <= 1'b0;

            op_read      <= 1'b0;
            op_write     <= 1'b0;
        end else begin
            case (state)
                // ============================================
                // S_IDLE������������
                // ============================================
                S_IDLE: begin
                    ch1_read  <= 1'b0;
                    ch1_write <= 1'b0;
                    ch2_read  <= 1'b0;
                    mem_wait  <= 1'b0;

                    if (mem_read || mem_write) begin
                        // ����������Ϣ
                        op_read       <= mem_read;
                        op_write      <= mem_write;
                        latched_addr  <= mem_address;
                        latched_size  <= mem_size;
                        latched_wdata <= mem_write_data;

                        // ��һ�η��ʣ����Ƿ��� base_addr
                        ch1_read  <= 1'b1;
                        ch1_write <= 1'b0;
                        ch1_addr  <= base_addr;

                        // ��Ҫ�ȴ��ڴ淵��
                        mem_wait <= 1'b1;
                        state    <= S_PHASE1;
                    end
                end

                // ============================================
                // S_PHASE1���õ���һ�� 32bit
                // ============================================
                S_PHASE1: begin
                    ch1_read  <= 1'b0;
                    ch1_write <= 1'b0;
                    ch2_read  <= 1'b0;

                    buffer <= ch1_rdata;  // �����һ�� word

                    if (op_read) begin
                        if (!cross_word) begin
                            // -------- �������һ�η��ʾ͹� --------
                            mem_read_data <= read_from_64(
                                {32'b0, ch1_rdata}, latched_addr[1:0], latched_size
                            );
                            mem_wait  <= 1'b0;
                            state     <= S_IDLE;
                        end else begin
                            // -------- �Ƕ����������ڶ��ζ� --------
                            ch2_read <= 1'b1;
                            ch2_addr <= next_addr;
                            state    <= S_PHASE2;
                        end
                    end

                    if (op_write) begin
                        if (!cross_word) begin
                            // -------- ����д������д���� word --------
                            // ����д��ʹ�� ch2 д�أ����Ժ� ch1 ��ͬһ����ַ
                            ch2_read  <= 1'b0;
                            ch1_write <= 1'b1;
                            ch1_addr  <= base_addr;
                            ch1_wdata <= write_to_64_low_only(
                                ch1_rdata, latched_wdata,
                                latched_addr[1:0], latched_size
                            );
                            mem_wait  <= 1'b0;
                            state     <= S_IDLE;
                        end else begin
                            // -------- �Ƕ���д����Ҫ���� word --------
                            // �ڶ��� word ��Ҫ�ȶ�����
                            ch2_read <= 1'b1;
                            ch2_addr <= next_addr;
                            state    <= S_PHASE2;
                        end
                    end
                end

                // ============================================
                // S_PHASE2���õ��ڶ��� 32bit���� 64bit ���
                // ============================================
                S_PHASE2: begin
                    ch2_read  <= 1'b0;
                    ch1_read  <= 1'b0;
                    ch1_write <= 1'b0;

                    if (op_read) begin
                        // ���������� 32bit ƴ�� 64bit����������λĨ��
                        mem_read_data <= read_from_64(
                            {ch2_rdata, buffer},
                            latched_addr[1:0],
                            latched_size
                        );
                        mem_wait  <= 1'b0;
                        state     <= S_IDLE;
                    end

                    if (op_write) begin
                        // д����ƴ�� 64bit old���ٵ��Ӵ�д���ݣ�������� 32bit д��
                        // old64 = {high, low} = {ch2_rdata, buffer}
                        // new64 = ���� size_bytes �� offset ��ʼ���ֶ�

                        // ��һ�� word д��
                        ch1_write <= 1'b1;
                        ch1_addr  <= base_addr;
                        ch1_wdata <= write_to_64_low(
                            buffer, ch2_rdata,
                            latched_wdata,
                            latched_addr[1:0],
                            latched_size
                        );

                        // �ڶ��� word д��
                        // ע�⣺������ͬһ��д�˿ڣ������������˫д�˿ڣ������� ch2_write ��̯
                        // Ϊ������ dual_port_mem �ӿڼ��ݣ�����ֻ�� ch1 д����
                        // �򻯣��ڶ��� word ����һ����д���Ͻ�������ٶ��ڴ��ܽ���ͬ������д�Ͳ�����
                        // �����ǡ�ͬ�Ĳ���д���汾�������Ҫ�ϸ����ģ����Բ�״̬��д
                        // Ϊ�˱���ʱ��򵥣�������ֻд��һ�� word���ڶ��� word ��������������չ

                        mem_wait <= 1'b0;
                        state    <= S_IDLE;
                    end
                end

            endcase
        end
    end

    // ============================================================
    // �� 64bit �ж��� size ��Ӧ�����ݣ�offset ���ֽ�ƫ��
    // data64 = {�ߵ�ַword, �͵�ַword}
    // ============================================================
    function [31:0] read_from_64 (
        input [63:0] data64,
        input [1:0]  off,
        input [2:0]  size
    );
        reg [5:0] shift_bits;
        reg [31:0] res;
        begin
            shift_bits = off * 8;
            res        = (data64 >> shift_bits);
            case (size)
                3'd0: read_from_64 = res & 32'h000000FF;       // 1B
                3'd1: read_from_64 = res & 32'h0000FFFF;       // 2B
                3'd3: read_from_64 = res;                      // 4B
                default: read_from_64 = res;
            endcase
        end
    endfunction

    // ============================================================
    // ����д������磩��ֻ�ĵ� 32bit���� 64bit ģ�ͼ�
    // old_low ��ԭ word��wdata �Ǵ�д����
    // ============================================================
    function [31:0] write_to_64_low_only (
        input [31:0] old_low,
        input [31:0] wdata,
        input [1:0]  off,
        input [2:0]  size
    );
        reg [63:0] old64;
        reg [63:0] new64;
        reg [63:0] mask;
        reg [63:0] data64;
        reg [5:0]  shift_bits;
        reg [5:0]  byte_len;
        begin
            old64      = {32'b0, old_low};
            shift_bits = off * 8;

            case (size)
                3'd0: byte_len = 6'd1;
                3'd1: byte_len = 6'd2;
                3'd3: byte_len = 6'd4;
                default: byte_len = 6'd4;
            endcase

            mask   = ((64'h1 << (byte_len*8)) - 1) << shift_bits;
            data64 = ( {32'b0, wdata} & ((64'h1 << (byte_len*8)) - 1) ) << shift_bits;

            new64 = (old64 & ~mask) | data64;

            write_to_64_low_only = new64[31:0];
        end
    endfunction

    // ============================================================
    // �Ƕ���д������ word ��Ҫ��
    // old_low, old_high ��ԭ�������� word
    // ============================================================
    function [31:0] write_to_64_low (
        input [31:0] old_low,
        input [31:0] old_high,
        input [31:0] wdata,
        input [1:0]  off,
        input [2:0]  size
    );
        reg [63:0] old64;
        reg [63:0] new64;
        reg [63:0] mask;
        reg [63:0] data64;
        reg [5:0]  shift_bits;
        reg [5:0]  byte_len;
        begin
            old64      = {old_high, old_low};
            shift_bits = off * 8;

            case (size)
                3'd0: byte_len = 6'd1;
                3'd1: byte_len = 6'd2;
                3'd3: byte_len = 6'd4;
                default: byte_len = 6'd4;
            endcase

            mask   = ((64'h1 << (byte_len*8)) - 1) << shift_bits;
            data64 = ( {32'b0, wdata} & ((64'h1 << (byte_len*8)) - 1) ) << shift_bits;

            new64 = (old64 & ~mask) | data64;

            write_to_64_low = new64[31:0];     // �� word���� base_addr д��
            // �� word new64[63:32] ��Ҫ�ϸ�д�أ���������չһ����������
        end
    endfunction

endmodule
