module ZXE6ZXA0ZX88z_2 (clk, rst, POP, PUSH, VALUE, OUTPUT);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] POP;
  input  wire [0:0] PUSH;
  input  wire [7:0] VALUE;
  output  wire [7:0] OUTPUT;

  TC_Switch # (.UUID(64'd4075459734019581736 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_0 (.en(wire_53), .in(wire_11), .out(OUTPUT));
  TC_Switch # (.UUID(64'd1743450744501712481 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_1 (.en(wire_1), .in(wire_118), .out(wire_30_1));
  TC_Nor # (.UUID(64'd2790480606642533264 ^ UUID), .BIT_WIDTH(64'd1)) Nor_2 (.in0(wire_53), .in1(wire_1), .out(wire_7));
  TC_Switch # (.UUID(64'd3620968006466173408 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_53), .in(wire_19), .out(wire_30_2));
  TC_Switch # (.UUID(64'd2715955857100762530 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_7), .in(wire_11), .out(wire_30_0));
  TC_Maker8 # (.UUID(64'd2469106912994579223 ^ UUID)) Maker8_5 (.in0(wire_37), .in1(wire_68), .in2(wire_25), .in3(wire_17), .in4(wire_57), .in5(wire_32), .in6(wire_61), .in7(wire_102), .out(wire_11));
  TC_Splitter8 # (.UUID(64'd127272120207574493 ^ UUID)) Splitter8_6 (.in(wire_30), .out0(wire_147), .out1(wire_127), .out2(wire_99), .out3(wire_139), .out4(wire_130), .out5(wire_41), .out6(wire_59), .out7(wire_39));
  TC_DelayLine # (.UUID(64'd3393656051382904683 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_7 (.clk(clk), .rst(rst), .in(wire_39), .out(wire_102));
  TC_DelayLine # (.UUID(64'd1334706193285872778 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_8 (.clk(clk), .rst(rst), .in(wire_59), .out(wire_61));
  TC_DelayLine # (.UUID(64'd1514987499206398818 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_9 (.clk(clk), .rst(rst), .in(wire_41), .out(wire_32));
  TC_DelayLine # (.UUID(64'd716467056116742491 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_10 (.clk(clk), .rst(rst), .in(wire_130), .out(wire_57));
  TC_DelayLine # (.UUID(64'd3104012118539659468 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_11 (.clk(clk), .rst(rst), .in(wire_139), .out(wire_17));
  TC_DelayLine # (.UUID(64'd3570369426499643292 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_12 (.clk(clk), .rst(rst), .in(wire_99), .out(wire_25));
  TC_DelayLine # (.UUID(64'd3526182291069794268 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_13 (.clk(clk), .rst(rst), .in(wire_127), .out(wire_68));
  TC_DelayLine # (.UUID(64'd1168041412397167956 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_14 (.clk(clk), .rst(rst), .in(wire_147), .out(wire_37));
  TC_DelayLine # (.UUID(64'd1205367239378628770 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_15 (.clk(clk), .rst(rst), .in(wire_92), .out(wire_70));
  TC_DelayLine # (.UUID(64'd3257161681445367497 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_16 (.clk(clk), .rst(rst), .in(wire_143), .out(wire_2));
  TC_DelayLine # (.UUID(64'd3574738129638164796 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_17 (.clk(clk), .rst(rst), .in(wire_58), .out(wire_10));
  TC_DelayLine # (.UUID(64'd3062098513855271243 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_18 (.clk(clk), .rst(rst), .in(wire_121), .out(wire_119));
  TC_DelayLine # (.UUID(64'd4405201251493582131 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_19 (.clk(clk), .rst(rst), .in(wire_134), .out(wire_80));
  TC_DelayLine # (.UUID(64'd4241083042292952884 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_20 (.clk(clk), .rst(rst), .in(wire_132), .out(wire_69));
  TC_DelayLine # (.UUID(64'd4510446554595175181 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_21 (.clk(clk), .rst(rst), .in(wire_111), .out(wire_89));
  TC_DelayLine # (.UUID(64'd591680535643659490 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_22 (.clk(clk), .rst(rst), .in(wire_43), .out(wire_135));
  TC_Splitter8 # (.UUID(64'd2141641741365277671 ^ UUID)) Splitter8_23 (.in(wire_15), .out0(wire_92), .out1(wire_143), .out2(wire_58), .out3(wire_121), .out4(wire_134), .out5(wire_132), .out6(wire_111), .out7(wire_43));
  TC_Maker8 # (.UUID(64'd772014627663534443 ^ UUID)) Maker8_24 (.in0(wire_70), .in1(wire_2), .in2(wire_10), .in3(wire_119), .in4(wire_80), .in5(wire_69), .in6(wire_89), .in7(wire_135), .out(wire_19));
  TC_Switch # (.UUID(64'd346468829949457959 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_1), .in(wire_11), .out(wire_15_1));
  TC_Switch # (.UUID(64'd1830357213095960909 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_7), .in(wire_19), .out(wire_15_0));
  TC_DelayLine # (.UUID(64'd248807222444607629 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_27 (.clk(clk), .rst(rst), .in(wire_122), .out(wire_123));
  TC_DelayLine # (.UUID(64'd802433610171549351 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_28 (.clk(clk), .rst(rst), .in(wire_56), .out(wire_22));
  TC_DelayLine # (.UUID(64'd3991703851828864956 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_105), .out(wire_141));
  TC_DelayLine # (.UUID(64'd4395842919601474748 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_30 (.clk(clk), .rst(rst), .in(wire_60), .out(wire_72));
  TC_DelayLine # (.UUID(64'd2005584888825114944 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_31 (.clk(clk), .rst(rst), .in(wire_125), .out(wire_38));
  TC_DelayLine # (.UUID(64'd2119628560784434773 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_32 (.clk(clk), .rst(rst), .in(wire_144), .out(wire_108));
  TC_DelayLine # (.UUID(64'd1850531147289421062 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_33 (.clk(clk), .rst(rst), .in(wire_5), .out(wire_83));
  TC_DelayLine # (.UUID(64'd4264777058425197048 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_34 (.clk(clk), .rst(rst), .in(wire_9), .out(wire_137));
  TC_Splitter8 # (.UUID(64'd1423284249291036898 ^ UUID)) Splitter8_35 (.in(wire_12), .out0(wire_122), .out1(wire_56), .out2(wire_105), .out3(wire_60), .out4(wire_125), .out5(wire_144), .out6(wire_5), .out7(wire_9));
  TC_Maker8 # (.UUID(64'd2472972256614238286 ^ UUID)) Maker8_36 (.in0(wire_123), .in1(wire_22), .in2(wire_141), .in3(wire_72), .in4(wire_38), .in5(wire_108), .in6(wire_83), .in7(wire_137), .out(wire_74));
  TC_Switch # (.UUID(64'd2996510639430170199 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_37 (.en(wire_1), .in(wire_19), .out(wire_12_0));
  TC_Switch # (.UUID(64'd3370806962555693786 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_38 (.en(wire_7), .in(wire_74), .out(wire_12_1));
  TC_DelayLine # (.UUID(64'd1482348844004579601 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_39 (.clk(clk), .rst(rst), .in(wire_104), .out(wire_117));
  TC_DelayLine # (.UUID(64'd2232322640709479327 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_40 (.clk(clk), .rst(rst), .in(wire_109), .out(wire_28));
  TC_DelayLine # (.UUID(64'd4068393948222517207 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_41 (.clk(clk), .rst(rst), .in(wire_120), .out(wire_100));
  TC_DelayLine # (.UUID(64'd3389451547221995772 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_42 (.clk(clk), .rst(rst), .in(wire_95), .out(wire_71));
  TC_DelayLine # (.UUID(64'd2734922808867655483 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_43 (.clk(clk), .rst(rst), .in(wire_145), .out(wire_20));
  TC_DelayLine # (.UUID(64'd3530346876910630963 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_44 (.clk(clk), .rst(rst), .in(wire_45), .out(wire_91));
  TC_DelayLine # (.UUID(64'd152115064831178903 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_45 (.clk(clk), .rst(rst), .in(wire_54), .out(wire_35));
  TC_DelayLine # (.UUID(64'd4282287041681468623 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_46 (.clk(clk), .rst(rst), .in(wire_88), .out(wire_136));
  TC_Splitter8 # (.UUID(64'd2996546740734991049 ^ UUID)) Splitter8_47 (.in(wire_31), .out0(wire_104), .out1(wire_109), .out2(wire_120), .out3(wire_95), .out4(wire_145), .out5(wire_45), .out6(wire_54), .out7(wire_88));
  TC_Maker8 # (.UUID(64'd2461916142859953651 ^ UUID)) Maker8_48 (.in0(wire_117), .in1(wire_28), .in2(wire_100), .in3(wire_71), .in4(wire_20), .in5(wire_91), .in6(wire_35), .in7(wire_136), .out(wire_49));
  TC_Switch # (.UUID(64'd3274850918193023928 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_1), .in(wire_74), .out(wire_31_1));
  TC_Switch # (.UUID(64'd3638538971750995833 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_7), .in(wire_49), .out(wire_31_0));
  TC_DelayLine # (.UUID(64'd78040464347862748 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_51 (.clk(clk), .rst(rst), .in(wire_0), .out(wire_76));
  TC_DelayLine # (.UUID(64'd2841552515341463628 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_52 (.clk(clk), .rst(rst), .in(wire_55), .out(wire_97));
  TC_DelayLine # (.UUID(64'd1573878953791415923 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_53 (.clk(clk), .rst(rst), .in(wire_112), .out(wire_106));
  TC_DelayLine # (.UUID(64'd1562778224091037259 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_54 (.clk(clk), .rst(rst), .in(wire_63), .out(wire_73));
  TC_DelayLine # (.UUID(64'd3173381059019276823 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_55 (.clk(clk), .rst(rst), .in(wire_128), .out(wire_33));
  TC_DelayLine # (.UUID(64'd2766581341910007777 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_56 (.clk(clk), .rst(rst), .in(wire_115), .out(wire_3));
  TC_DelayLine # (.UUID(64'd3338101237389752377 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_57 (.clk(clk), .rst(rst), .in(wire_8), .out(wire_142));
  TC_DelayLine # (.UUID(64'd1987811693578649385 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_58 (.clk(clk), .rst(rst), .in(wire_85), .out(wire_21));
  TC_Splitter8 # (.UUID(64'd4524465079344680757 ^ UUID)) Splitter8_59 (.in(wire_16), .out0(wire_0), .out1(wire_55), .out2(wire_112), .out3(wire_63), .out4(wire_128), .out5(wire_115), .out6(wire_8), .out7(wire_85));
  TC_Maker8 # (.UUID(64'd2966218995392052499 ^ UUID)) Maker8_60 (.in0(wire_76), .in1(wire_97), .in2(wire_106), .in3(wire_73), .in4(wire_33), .in5(wire_3), .in6(wire_142), .in7(wire_21), .out(wire_51));
  TC_Switch # (.UUID(64'd3754574919523500658 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_61 (.en(wire_1), .in(wire_49), .out(wire_16_0));
  TC_Switch # (.UUID(64'd4079238810151005972 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_62 (.en(wire_7), .in(wire_51), .out(wire_16_2));
  TC_DelayLine # (.UUID(64'd2781728321311578945 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_63 (.clk(clk), .rst(rst), .in(wire_101), .out(wire_65));
  TC_DelayLine # (.UUID(64'd1631081794559958622 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_64 (.clk(clk), .rst(rst), .in(wire_14), .out(wire_98));
  TC_DelayLine # (.UUID(64'd2403130787508255652 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_65 (.clk(clk), .rst(rst), .in(wire_48), .out(wire_124));
  TC_DelayLine # (.UUID(64'd1663662469583701893 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_66 (.clk(clk), .rst(rst), .in(wire_86), .out(wire_107));
  TC_DelayLine # (.UUID(64'd2001633194596840400 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_67 (.clk(clk), .rst(rst), .in(wire_146), .out(wire_133));
  TC_DelayLine # (.UUID(64'd3987881675664836630 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_68 (.clk(clk), .rst(rst), .in(wire_26), .out(wire_40));
  TC_DelayLine # (.UUID(64'd1278355622528026551 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_69 (.clk(clk), .rst(rst), .in(wire_126), .out(wire_79));
  TC_DelayLine # (.UUID(64'd4117982776272952303 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_70 (.clk(clk), .rst(rst), .in(wire_66), .out(wire_110));
  TC_Splitter8 # (.UUID(64'd4571229142849269409 ^ UUID)) Splitter8_71 (.in(wire_23), .out0(wire_101), .out1(wire_14), .out2(wire_48), .out3(wire_86), .out4(wire_146), .out5(wire_26), .out6(wire_126), .out7(wire_66));
  TC_Maker8 # (.UUID(64'd2150865959364266972 ^ UUID)) Maker8_72 (.in0(wire_65), .in1(wire_98), .in2(wire_124), .in3(wire_107), .in4(wire_133), .in5(wire_40), .in6(wire_79), .in7(wire_110), .out(wire_4));
  TC_Switch # (.UUID(64'd2665755057558486683 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_73 (.en(wire_1), .in(wire_51), .out(wire_23_1));
  TC_Switch # (.UUID(64'd2597763441492845171 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_74 (.en(wire_7), .in(wire_4), .out(wire_23_0));
  TC_DelayLine # (.UUID(64'd3967024153069262303 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_75 (.clk(clk), .rst(rst), .in(wire_29), .out(wire_84));
  TC_DelayLine # (.UUID(64'd972683716322260849 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_76 (.clk(clk), .rst(rst), .in(wire_103), .out(wire_140));
  TC_DelayLine # (.UUID(64'd1986549943731871725 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_77 (.clk(clk), .rst(rst), .in(wire_87), .out(wire_62));
  TC_DelayLine # (.UUID(64'd2630879542408606380 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_78 (.clk(clk), .rst(rst), .in(wire_6), .out(wire_24));
  TC_DelayLine # (.UUID(64'd857310293201125423 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_79 (.clk(clk), .rst(rst), .in(wire_116), .out(wire_47));
  TC_DelayLine # (.UUID(64'd1664653121859202556 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_80 (.clk(clk), .rst(rst), .in(wire_18), .out(wire_77));
  TC_DelayLine # (.UUID(64'd1277125745797389229 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_81 (.clk(clk), .rst(rst), .in(wire_131), .out(wire_81));
  TC_DelayLine # (.UUID(64'd1974208262777888759 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_82 (.clk(clk), .rst(rst), .in(wire_93), .out(wire_138));
  TC_Splitter8 # (.UUID(64'd2449185560105409524 ^ UUID)) Splitter8_83 (.in(wire_36), .out0(wire_29), .out1(wire_103), .out2(wire_87), .out3(wire_6), .out4(wire_116), .out5(wire_18), .out6(wire_131), .out7(wire_93));
  TC_Maker8 # (.UUID(64'd2540742893926616621 ^ UUID)) Maker8_84 (.in0(wire_84), .in1(wire_140), .in2(wire_62), .in3(wire_24), .in4(wire_47), .in5(wire_77), .in6(wire_81), .in7(wire_138), .out(wire_46));
  TC_Switch # (.UUID(64'd4237025915478602165 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_85 (.en(wire_1), .in(wire_4), .out(wire_36_1));
  TC_Switch # (.UUID(64'd3757407907371428479 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_86 (.en(wire_7), .in(wire_46), .out(wire_36_0));
  TC_DelayLine # (.UUID(64'd251654647185254920 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_87 (.clk(clk), .rst(rst), .in(wire_82), .out(wire_13));
  TC_DelayLine # (.UUID(64'd1903788780711488873 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_88 (.clk(clk), .rst(rst), .in(wire_64), .out(wire_113));
  TC_DelayLine # (.UUID(64'd1820407957447023659 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_89 (.clk(clk), .rst(rst), .in(wire_44), .out(wire_42));
  TC_DelayLine # (.UUID(64'd4133323914555002002 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_90 (.clk(clk), .rst(rst), .in(wire_94), .out(wire_50));
  TC_DelayLine # (.UUID(64'd3804304960686378029 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_91 (.clk(clk), .rst(rst), .in(wire_96), .out(wire_67));
  TC_DelayLine # (.UUID(64'd493552682330002982 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_92 (.clk(clk), .rst(rst), .in(wire_75), .out(wire_27));
  TC_DelayLine # (.UUID(64'd1957394206760702121 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_93 (.clk(clk), .rst(rst), .in(wire_129), .out(wire_114));
  TC_DelayLine # (.UUID(64'd1626460170447878873 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_94 (.clk(clk), .rst(rst), .in(wire_52), .out(wire_78));
  TC_Splitter8 # (.UUID(64'd200448370920329985 ^ UUID)) Splitter8_95 (.in(wire_90), .out0(wire_82), .out1(wire_64), .out2(wire_44), .out3(wire_94), .out4(wire_96), .out5(wire_75), .out6(wire_129), .out7(wire_52));
  TC_Maker8 # (.UUID(64'd3193589546896296758 ^ UUID)) Maker8_96 (.in0(wire_13), .in1(wire_113), .in2(wire_42), .in3(wire_50), .in4(wire_67), .in5(wire_27), .in6(wire_114), .in7(wire_78), .out(wire_34));
  TC_Switch # (.UUID(64'd1122850571013921338 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_97 (.en(wire_1), .in(wire_46), .out(wire_90_0));
  TC_Switch # (.UUID(64'd3170085125241982752 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_98 (.en(wire_7), .in(wire_34), .out(wire_90_1));
  TC_Switch # (.UUID(64'd3971553172260668966 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_99 (.en(wire_53), .in(wire_74), .out(wire_15_2));
  TC_Switch # (.UUID(64'd3069202300250339585 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_100 (.en(wire_53), .in(wire_49), .out(wire_12_2));
  TC_Switch # (.UUID(64'd2675741184577763658 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_101 (.en(wire_53), .in(wire_51), .out(wire_31_2));
  TC_Switch # (.UUID(64'd1824493707107369539 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_102 (.en(wire_53), .in(wire_4), .out(wire_16_1));
  TC_Switch # (.UUID(64'd2159838870751308370 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_103 (.en(wire_53), .in(wire_46), .out(wire_23_2));
  TC_Switch # (.UUID(64'd3883996631719742858 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_104 (.en(wire_53), .in(wire_34), .out(wire_36_2));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  assign wire_1 = PUSH;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_12_0;
  wire [7:0] wire_12_1;
  wire [7:0] wire_12_2;
  assign wire_12 = wire_12_0|wire_12_1|wire_12_2;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_15_0;
  wire [7:0] wire_15_1;
  wire [7:0] wire_15_2;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2;
  wire [7:0] wire_16;
  wire [7:0] wire_16_0;
  wire [7:0] wire_16_1;
  wire [7:0] wire_16_2;
  assign wire_16 = wire_16_0|wire_16_1|wire_16_2;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_23_0;
  wire [7:0] wire_23_1;
  wire [7:0] wire_23_2;
  assign wire_23 = wire_23_0|wire_23_1|wire_23_2;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_30_0;
  wire [7:0] wire_30_1;
  wire [7:0] wire_30_2;
  assign wire_30 = wire_30_0|wire_30_1|wire_30_2;
  wire [7:0] wire_31;
  wire [7:0] wire_31_0;
  wire [7:0] wire_31_1;
  wire [7:0] wire_31_2;
  assign wire_31 = wire_31_0|wire_31_1|wire_31_2;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [7:0] wire_36_0;
  wire [7:0] wire_36_1;
  wire [7:0] wire_36_2;
  assign wire_36 = wire_36_0|wire_36_1|wire_36_2;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [7:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  assign wire_53 = POP;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [7:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [7:0] wire_90;
  wire [7:0] wire_90_0;
  wire [7:0] wire_90_1;
  assign wire_90 = wire_90_0|wire_90_1;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [7:0] wire_118;
  assign wire_118 = VALUE;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [0:0] wire_126;
  wire [0:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [0:0] wire_131;
  wire [0:0] wire_132;
  wire [0:0] wire_133;
  wire [0:0] wire_134;
  wire [0:0] wire_135;
  wire [0:0] wire_136;
  wire [0:0] wire_137;
  wire [0:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [0:0] wire_141;
  wire [0:0] wire_142;
  wire [0:0] wire_143;
  wire [0:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [0:0] wire_147;

endmodule
